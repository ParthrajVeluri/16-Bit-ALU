Library ieee; 
Use ieee.std_logic_1164.all;

Entity latch1 is 
	Port (A: in std_logic_vector(7 downto 0);
			Resetn,Clock: in std_logic;
			Q : out std_logic_vector(7 downto 0));
end latch1; 

Architecture Behaviour of latch1 is 
Begin 
	Process (Resetn, Clock)
	Begin 
		If Resetn = '0' then 
			Q <= "00000000";
		elsif Clock'EVENT AND Clock = '1' then 
			Q <= A; 
		end if; 
	end process; 
end Behaviour;
